axi_bfm.sv
module_axi_slave.sv
axi_tb_top.sv
