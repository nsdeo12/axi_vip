`include "axi_slave.sv"
`include "byte_tx.sv"
`include "axi_if.sv"
`include "axi_transaction.sv"
`include "axi_tx_resp.sv"
`include "axi_monitor.sv"
//`include "axi_ref.sv"
//`include "axi_cov.sv"
`include "axi_bfm.sv"
`include "axi_gen.sv"
`include "axi_env.sv"
`include "axi_tb.sv"
`include "axi_tb_top.sv"
