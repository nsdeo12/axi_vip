class axi_ckr;

endclass
